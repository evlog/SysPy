----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:13:13 10/22/2011 
-- Design Name: 
-- Module Name:    datamemddr5forLEON - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity datamemddr5forLEON is
port (clk : in std_logic; 
 	--we  : in std_logic; 
 	en,restart,enfroFSM,sendnext  : in std_logic;
 	ce2int : out std_logic;
	muxgpio: out std_logic_vector(1 downto 0);
	di2,dii2,dii3,dii4   : in std_logic_vector(15 downto 0);
 	--a: in std_logic_vector(8 downto 0); 
 	di,dii,diii,diiii  : in std_logic_vector(287 downto 0); 
	doid,dooid,doooid,dooooid:out std_logic_vector(8 downto 0);
 	do,do0,do1,do2,do3,do4,do5,do6,do7,doo,doo0,doo1,doo2,doo3,doo4,doo5,doo6,doo7,dooo,dooo0,dooo1,dooo2,dooo3,dooo4,dooo5,dooo6,dooo7,doooo,doooo0,doooo1,doooo2,doooo3,doooo4,doooo5,doooo6,doooo7  : out std_logic_vector(31 downto 0));
end datamemddr5forLEON;

architecture Behavioral of datamemddr5forLEON is

signal we,we2,we3,we4 : std_logic:='0';
signal acnt,acnt2,acnt3,acnt4:std_logic_vector(8 downto 0):="000000000";
--type states is(s_delay,s_update1,s_update2,s_update1a,s_update2a,s_update1b,s_update2b,s_update1c,s_update2c,s_started,s_starteda,s_begin1,s_start1,s_start2a,s_start2,s_start3,s_start4a,s_start4,s_start5,s_start6a,s_start6,s_start7,s_start8a,s_start8,s_1, s_2, s_3,s_4,s_5,s_6,s_7,s_8,s_9,s_10);
type states is(s_start0,s_start1,s_start2,s_start3,s_start4a,s_start4,s_start5,s_start6a,s_start6,s_start7,s_start8a,s_start8,s_start9,s_start10,s_start11,s_start12,s_start13,s_start14,s_start15,s_start16,s_start17,s_start18,s_start19,s_start20,s_start21,s_start22,s_start23,s_start24,s_start25,s_start26,s_start27,s_start28,s_start29,s_start30,s_start31,s_start32);
signal state, previous_state: states;

type ram_type is array(0 to 511) of std_logic_vector(287 downto 0);
signal RAM:ram_type:=
(X"0000000a00000012000000123A83126E0000000300000012000000120000001200000012", X"00000003000000120000001238D1B7170000000900000012000000120000001200000012", X"0000000200000012000000123A01C2E300000002000000110000000e0000001200000012", X"00000000000000120000001238D1B7170000000000000002000000100000001200000012", X"00000006000000120000001238D1B7170000000600000002000000100000001200000012", X"00000002000000120000001238D1B717000000090000000f000000120000001200000012",X"00000011000000120000001239E30446000000090000000d000000120000001200000012", X"0000000300000012000000123BC49BA500000000000000030000000c0000001200000012", X"0000000100000012000000123A5844D0000000110000000b000000120000001200000012", X"0000000000000011000000123A97635E0000000100000012000000120000001200000012",  
 X"0000000100000012000000123741C6DF0000000000000011000000120000001200000012", X"0000001200000012000000123DA3D70A0000000800000012000000120000001200000012", X"00000008000000120000001237A7C5AC0000000900000013000000120000001200000012", X"00000008000000050000001238D1B7170000000800000004000000120000001200000012", X"0000000000000004000000123A03126E0000000600000004000000120000001200000012", X"0000000600000012000000123f0000000000000000000012000000120000001200000012",X"000000110000000400000012400000000000000700000004000000120000001200000012", X"0000000700000012000000123f0000000000001100000012000000120000001200000012", X"00000007000000120000001239E30446000000090000000d000000120000001200000012", X"0000000400000012000000123A03126E0000000500000012000000120000001200000012",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001");

type ram_type2 is array(0 to 511) of std_logic_vector(15 downto 0);
signal RAM2:ram_type2:= 
(X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008");
 
 type ram_type3 is array(0 to 511) of std_logic_vector(287 downto 0);
signal RAM3:ram_type3:=
(X"0000000a00000012000000123A83126E0000000300000012000000120000001200000012", X"00000003000000120000001238D1B7170000000900000012000000120000001200000012", X"0000000200000012000000123A01C2E300000002000000110000000e0000001200000012", X"00000000000000120000001238D1B7170000000000000002000000100000001200000012", X"00000006000000120000001238D1B7170000000600000002000000100000001200000012", X"00000002000000120000001238D1B717000000090000000f000000120000001200000012",X"00000011000000120000001239E30446000000090000000d000000120000001200000012", X"0000000300000012000000123BC49BA500000000000000030000000c0000001200000012", X"0000000100000012000000123A5844D0000000110000000b000000120000001200000012", X"0000000000000011000000123A97635E0000000100000012000000120000001200000012",  
 X"0000000100000012000000123741C6DF0000000000000011000000120000001200000012", X"0000001200000012000000123DA3D70A0000000800000012000000120000001200000012", X"00000008000000120000001237A7C5AC0000000900000013000000120000001200000012", X"00000008000000050000001238D1B7170000000800000004000000120000001200000012", X"0000000000000004000000123A03126E0000000600000004000000120000001200000012", X"0000000600000012000000123f0000000000000000000012000000120000001200000012",X"000000110000000400000012400000000000000700000004000000120000001200000012", X"0000000700000012000000123f0000000000001100000012000000120000001200000012", X"00000007000000120000001239E30446000000090000000d000000120000001200000012", X"0000000400000012000000123A03126E0000000500000012000000120000001200000012",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001");

type ram_type4 is array(0 to 511) of std_logic_vector(15 downto 0);
signal RAM4:ram_type4:= 
(X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008");
 
type ram_type5 is array(0 to 511) of std_logic_vector(287 downto 0);
signal RAM5:ram_type5:=
(X"0000000a00000012000000123A83126E0000000300000012000000120000001200000012", X"00000003000000120000001238D1B7170000000900000012000000120000001200000012", X"0000000200000012000000123A01C2E300000002000000110000000e0000001200000012", X"00000000000000120000001238D1B7170000000000000002000000100000001200000012", X"00000006000000120000001238D1B7170000000600000002000000100000001200000012", X"00000002000000120000001238D1B717000000090000000f000000120000001200000012",X"00000011000000120000001239E30446000000090000000d000000120000001200000012", X"0000000300000012000000123BC49BA500000000000000030000000c0000001200000012", X"0000000100000012000000123A5844D0000000110000000b000000120000001200000012", X"0000000000000011000000123A97635E0000000100000012000000120000001200000012",  
 X"0000000100000012000000123741C6DF0000000000000011000000120000001200000012", X"0000001200000012000000123DA3D70A0000000800000012000000120000001200000012", X"00000008000000120000001237A7C5AC0000000900000013000000120000001200000012", X"00000008000000050000001238D1B7170000000800000004000000120000001200000012", X"0000000000000004000000123A03126E0000000600000004000000120000001200000012", X"0000000600000012000000123f0000000000000000000012000000120000001200000012",X"000000110000000400000012400000000000000700000004000000120000001200000012", X"0000000700000012000000123f0000000000001100000012000000120000001200000012", X"00000007000000120000001239E30446000000090000000d000000120000001200000012", X"0000000400000012000000123A03126E0000000500000012000000120000001200000012",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001");

type ram_type6 is array(0 to 511) of std_logic_vector(15 downto 0);
signal RAM6:ram_type6:= 
(X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008");

type ram_type7 is array(0 to 511) of std_logic_vector(287 downto 0);
signal RAM7:ram_type7:=
(X"0000000a00000012000000123A83126E0000000300000012000000120000001200000012", X"00000003000000120000001238D1B7170000000900000012000000120000001200000012", X"0000000200000012000000123A01C2E300000002000000110000000e0000001200000012", X"00000000000000120000001238D1B7170000000000000002000000100000001200000012", X"00000006000000120000001238D1B7170000000600000002000000100000001200000012", X"00000002000000120000001238D1B717000000090000000f000000120000001200000012",X"00000011000000120000001239E30446000000090000000d000000120000001200000012", X"0000000300000012000000123BC49BA500000000000000030000000c0000001200000012", X"0000000100000012000000123A5844D0000000110000000b000000120000001200000012", X"0000000000000011000000123A97635E0000000100000012000000120000001200000012",  
 X"0000000100000012000000123741C6DF0000000000000011000000120000001200000012", X"0000001200000012000000123DA3D70A0000000800000012000000120000001200000012", X"00000008000000120000001237A7C5AC0000000900000013000000120000001200000012", X"00000008000000050000001238D1B7170000000800000004000000120000001200000012", X"0000000000000004000000123A03126E0000000600000004000000120000001200000012", X"0000000600000012000000123f0000000000000000000012000000120000001200000012",X"000000110000000400000012400000000000000700000004000000120000001200000012", X"0000000700000012000000123f0000000000001100000012000000120000001200000012", X"00000007000000120000001239E30446000000090000000d000000120000001200000012", X"0000000400000012000000123A03126E0000000500000012000000120000001200000012",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001");

type ram_type8 is array(0 to 511) of std_logic_vector(15 downto 0);
signal RAM8:ram_type8:= 
(X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008");
 
 type ram_type9 is array(0 to 511) of std_logic_vector(287 downto 0);
signal RAM9:ram_type9:=
(X"0000000a00000012000000123A83126E0000000300000012000000120000001200000012", X"00000003000000120000001238D1B7170000000900000012000000120000001200000012", X"0000000200000012000000123A01C2E300000002000000110000000e0000001200000012", X"00000000000000120000001238D1B7170000000000000002000000100000001200000012", X"00000006000000120000001238D1B7170000000600000002000000100000001200000012", X"00000002000000120000001238D1B717000000090000000f000000120000001200000012",X"00000011000000120000001239E30446000000090000000d000000120000001200000012", X"0000000300000012000000123BC49BA500000000000000030000000c0000001200000012", X"0000000100000012000000123A5844D0000000110000000b000000120000001200000012", X"0000000000000011000000123A97635E0000000100000012000000120000001200000012",  
 X"0000000100000012000000123741C6DF0000000000000011000000120000001200000012", X"0000001200000012000000123DA3D70A0000000800000012000000120000001200000012", X"00000008000000120000001237A7C5AC0000000900000013000000120000001200000012", X"00000008000000050000001238D1B7170000000800000004000000120000001200000012", X"0000000000000004000000123A03126E0000000600000004000000120000001200000012", X"0000000600000012000000123f0000000000000000000012000000120000001200000012",X"000000110000000400000012400000000000000700000004000000120000001200000012", X"0000000700000012000000123f0000000000001100000012000000120000001200000012", X"00000007000000120000001239E30446000000090000000d000000120000001200000012", X"0000000400000012000000123A03126E0000000500000012000000120000001200000012",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001");

type ram_type10 is array(0 to 511) of std_logic_vector(15 downto 0);
signal RAM10:ram_type10:= 
(X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008", 
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",  
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008", X"0008", X"0008", X"0008", X"0008",X"0008",X"0008", X"0008", X"0008",
 X"0008", X"0008");

begin 
process(clk,acnt,restart,enfroFSM)
 begin
  if clk'event and clk='1' then
  
    case state is
	 
	 when s_start0=>
	  ce2int<='0';muxgpio<="00";
   if acnt="111111111" then
	   acnt<="000000000";acnt2<="000000000";acnt3<="000000000";acnt4<="000000000";
	   state<=s_start1;
	 else
	 if enfroFSM='1' then
	  we <= '1';we2<='1';we3<='1';we4<='1';
     acnt<=acnt+1;acnt2<=acnt2+1;acnt3<=acnt3+1;acnt4<=acnt4+1;
	  else
	   we <= '0';we2<='0';we3<='0';we4<='0';
     acnt<=acnt;acnt2<=acnt2;acnt3<=acnt3;acnt4<=acnt4;
     end if;
     state<=s_start0;
	 end if; 
	  
	  when s_start1=>
	  ce2int<='1';muxgpio<="00";
   if acnt2="111111111" then
	   acnt<="000000000";acnt2<="000000000";acnt3<="000000000";acnt4<="000000000";
	   if restart='1' then
	   state<=s_start0;
	   else
       state<=s_start2;
      end if;
	 else
	  we <= '0';we3<='0';we4<='0';
	  if sendnext='1' then
     acnt<=acnt+1;
	  else
	  acnt<=acnt;acnt3<=acnt3;acnt4<=acnt4;
	  end if;
	  if enfroFSM='1' then
	  we2 <= '1';
     acnt2<=acnt2+1;
	  else
	   we2<='0';
      acnt2<=acnt2;
     end if;
     state<=s_start1;
	end if;
	
	when s_start2=>
	  ce2int<='1';muxgpio<="01";
   if acnt3="111111111" then
	   acnt<="000000000";acnt2<="000000000";acnt3<="000000000";acnt4<="000000000";
	   if restart='1' then
	   state<=s_start0;
	   else
       state<=s_start3;
      end if;
	 else
	  we2 <= '0';
	  if sendnext='1' then
     acnt2<=acnt2+1;
	  else
	  acnt2<=acnt2;
	  end if;
	  if enfroFSM='1' then
	  we3 <= '1';
     acnt3<=acnt3+1;
	  else
	   we3<='0';
      acnt3<=acnt3;
     end if;
     state<=s_start2;
	end if;
	
	when s_start3=>
	  ce2int<='1';muxgpio<="10";
   if acnt4="111111111" then
	   acnt<="000000000";acnt2<="000000000";acnt3<="000000000";acnt4<="000000000";
	   if restart='1' then
	   state<=s_start0;
	   else
       state<=s_start4;
      end if;
	 else
	  we3 <= '0';
	  if sendnext='1' then
     acnt3<=acnt3+1;
	  else
	  acnt3<=acnt3;
	  end if;
	  if enfroFSM='1' then
	  we4 <= '1';
     acnt4<=acnt4+1;
	  else
	   we4<='0';
      acnt4<=acnt4;
     end if;
     state<=s_start3;
	end if;
	
	when s_start4=>
	  ce2int<='1';muxgpio<="11";
   if acnt="111111111" then
	   acnt<="000000000";acnt2<="000000000";acnt3<="000000000";acnt4<="000000000";
	   if restart='1' then
	   state<=s_start0;
	   else
       state<=s_start1;
      end if;
	 else
	  we4 <= '0';
	  if sendnext='1' then
     acnt4<=acnt4+1;
	  else
	  acnt4<=acnt4;
	  end if;
	  if enfroFSM='1' then
	  we <= '1';
     acnt<=acnt+1;
	  else
	   we<='0';
      acnt<=acnt;
     end if;
     state<=s_start4;
	end if;
     	 
	  when others =>
        state<=s_start0;
		 
	end case;
	 
   end if;
end process;	


A1: process (clk,en,we) 
 begin 
if en='1' then
  if (clk'event and clk = '1') then
 	  --if en='1' then
 	   	if (we = '1') then 
 			RAM(conv_integer(acnt)) <= di; 
			RAM2(conv_integer(acnt)) <= di2;
 		else
		    do(31 downto 0)  <= RAM(conv_integer(acnt))(287 downto 256);
			 do0(31 downto 0) <= RAM(conv_integer(acnt))(255 downto 224);
		    do1(31 downto 0) <= RAM(conv_integer(acnt))(223 downto 192);
		    do2(31 downto 0) <= RAM(conv_integer(acnt))(191 downto 160);
 			 do3(31 downto 0) <= RAM(conv_integer(acnt))(159 downto 128);
			 do4(31 downto 0) <= RAM(conv_integer(acnt))(127 downto 96);
			 do5(31 downto 0) <= RAM(conv_integer(acnt))(95 downto 64);
			 do6(31 downto 0) <= RAM(conv_integer(acnt))(63 downto 32);
			 do7(31 downto 0) <= RAM(conv_integer(acnt))(31 downto 0);
			 doid<= RAM2(conv_integer(acnt))(8 downto 0);
 		end if;	  
 	end if; 
  end if;	
 end process; 
 
A2: process (clk,en,we2) 
 begin 
if en='1' then
  if (clk'event and clk = '1') then
 	  --if en='1' then
 	   	if (we2 = '1') then 
 			RAM3(conv_integer(acnt2)) <= dii; 
			RAM4(conv_integer(acnt2)) <= dii2;
 		else
		    doo(31 downto 0)  <= RAM3(conv_integer(acnt2))(287 downto 256);
			 doo0(31 downto 0) <= RAM3(conv_integer(acnt2))(255 downto 224);
		    doo1(31 downto 0) <= RAM3(conv_integer(acnt2))(223 downto 192);
		    doo2(31 downto 0) <= RAM3(conv_integer(acnt2))(191 downto 160);
 			 doo3(31 downto 0) <= RAM3(conv_integer(acnt2))(159 downto 128);
			 doo4(31 downto 0) <= RAM3(conv_integer(acnt2))(127 downto 96);
			 doo5(31 downto 0) <= RAM3(conv_integer(acnt2))(95 downto 64);
			 doo6(31 downto 0) <= RAM3(conv_integer(acnt2))(63 downto 32);
			 doo7(31 downto 0) <= RAM3(conv_integer(acnt2))(31 downto 0);
			 dooid<= RAM4(conv_integer(acnt2))(8 downto 0);
 		end if;	  
 	end if; 
  end if;	
 end process; 
 
 A3: process (clk,en,we3) 
 begin 
if en='1' then
  if (clk'event and clk = '1') then
 	  --if en='1' then
 	   	if (we3= '1') then 
 			RAM5(conv_integer(acnt3)) <= diii; 
			RAM6(conv_integer(acnt3)) <= dii3;
 		else
		    dooo(31 downto 0)  <= RAM5(conv_integer(acnt3))(287 downto 256);
			 dooo0(31 downto 0) <= RAM5(conv_integer(acnt3))(255 downto 224);
		    dooo1(31 downto 0) <= RAM5(conv_integer(acnt3))(223 downto 192);
		    dooo2(31 downto 0) <= RAM5(conv_integer(acnt3))(191 downto 160);
 			 dooo3(31 downto 0) <= RAM5(conv_integer(acnt3))(159 downto 128);
			 dooo4(31 downto 0) <= RAM5(conv_integer(acnt3))(127 downto 96);
			 dooo5(31 downto 0) <= RAM5(conv_integer(acnt3))(95 downto 64);
			 dooo6(31 downto 0) <= RAM5(conv_integer(acnt3))(63 downto 32);
			 dooo7(31 downto 0) <= RAM5(conv_integer(acnt3))(31 downto 0);
			 doooid<= RAM6(conv_integer(acnt3))(8 downto 0);
 		end if;	  
 	end if; 
  end if;	
 end process; 
 
 A4: process (clk,en,we4) 
 begin 
if en='1' then
  if (clk'event and clk = '1') then
 	  --if en='1' then
 	   	if (we4= '1') then 
 			RAM7(conv_integer(acnt4)) <= diiii; 
			RAM8(conv_integer(acnt4)) <= dii4;
 		else
		    doooo(31 downto 0)  <= RAM7(conv_integer(acnt4))(287 downto 256);
			 doooo0(31 downto 0) <= RAM7(conv_integer(acnt4))(255 downto 224);
		    doooo1(31 downto 0) <= RAM7(conv_integer(acnt4))(223 downto 192);
		    doooo2(31 downto 0) <= RAM7(conv_integer(acnt4))(191 downto 160);
 			 doooo3(31 downto 0) <= RAM7(conv_integer(acnt4))(159 downto 128);
			 doooo4(31 downto 0) <= RAM7(conv_integer(acnt4))(127 downto 96);
			 doooo5(31 downto 0) <= RAM7(conv_integer(acnt4))(95 downto 64);
			 doooo6(31 downto 0) <= RAM7(conv_integer(acnt4))(63 downto 32);
			 doooo7(31 downto 0) <= RAM7(conv_integer(acnt4))(31 downto 0);
			 dooooid<= RAM8(conv_integer(acnt4))(8 downto 0);
 		end if;	  
 	end if; 
  end if;	
 end process; 

end Behavioral;

