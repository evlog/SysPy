/home/SysPy_test/SysPy_ver/Python_script/paramsocs/LEONGILL/Addrepeatedly.vhd