----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    03:01:39 04/21/2011 
-- Design Name: 
-- Module Name:    Initmems - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Initmems is
port (clk : in std_logic; 
 	we  : in std_logic;
 	a   : in std_logic_vector(8 downto 0); 
 	di  : in std_logic_vector (159 downto 0); 
 	do  : out std_logic_vector(159 downto 0));
end Initmems;

architecture Behavioral of Initmems is
type ram_type is array(0 to 511) of std_logic_vector(159 downto 0);
signal RAM:ram_type:=
(X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e",
 X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a",X"00000001000000323E4CCCCC0000000B0000001e", X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a", X"00000001000000323E4CCCCC0000000B0000001e", 
 X"00000005000000643C23D70A000000160000003c", X"00000009000000963B83126E000000210000005a");
begin
process(clk,we)
begin
 if clk'event and clk='1' then
   if we='1' then
	  RAM(conv_integer(a))<=di;
	 else
     do<= RAM(conv_integer(a));	 
	end if;  
end if;
end process;	

end Behavioral;

