----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    07:25:44 09/14/2011 
-- Design Name: 
-- Module Name:    RTBIOMODEL189 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity RTBIOMODEL189 is
port (clk : in std_logic; 
 	we  : in std_logic; 
 	en  : in std_logic;
 	--ssr : in std_logic;
 	a   : in std_logic_vector(8 downto 0); 
 	di  : in std_logic_vector(287 downto 0); 
 	do,do0,do1,do2,do3,do4,do5,do6,do7  : out std_logic_vector(31 downto 0));
end RTBIOMODEL189;

architecture Behavioral of RTBIOMODEL189 is

type ram_type is array(0 to 511) of std_logic_vector(287 downto 0);
signal RAM:ram_type:=
(X"0000000300000012000000123A01C2E300000003000000000000000c0000001200000012", X"00000001000000120000001238D1B71700000001000000030000000e0000001200000012", X"00000003000000120000001238D1B717000000070000000d000000120000001200000012", X"00000000000000120000001239E30446000000070000000b000000120000001200000012", X"0000000800000012000000123D9FBE76000000010000000a000000120000001200000012", X"0000000200000012000000123A5844D00000000000000009000000120000001200000012",X"0000000100000000000000123A97635E0000000200000012000000120000001200000012", X"00000002000000120000001238F238970000000100000000000000120000001200000012", X"0000001200000012000000123DA3D70A000000060000000f000000120000001200000012", X"0000000600000012000000123851B7170000000700000012000000120000001200000012",  
 X"000000060000001200000012380A697A0000000600000004000000120000001200000012", X"0000000400000000000000123C23D70A0000000500000012000000120000001200000012", X"0000000500000012000000123A83126E000000040000000b000000120000001200000012", X"00000004000000120000001238D1B7170000000700000012000000120000001200000012", X"000000120000001200000012000000000000001200000012000000120000001200000012", X"000000120000001200000012000000000000001200000012000000120000001200000012",X"0000000900000089000000893189705F0000000800000081000000890000008900000089", X"0000008100000008000000893009705F0000000900000089000000890000008900000089", X"00000009000000890000008937A7C5AC0000000900000063000000890000008900000089", X"0000000a000000890000008931CE288E0000000900000081000000890000008900000089",
 X"0000008100000009000000893009705F0000000a00000089000000890000008900000089", X"0000000a000000890000008937A7C5AC0000000a00000063000000890000008900000089", X"0000000b00000089000000893189705F0000000a00000081000000890000008900000089", X"000000810000000a000000893009705F0000000b00000089000000890000008900000089", X"0000000b000000890000008937A7C5AC0000000b00000063000000890000008900000089", X"0000000c000000890000008931CE288E0000000b00000081000000890000008900000089",X"000000810000000b000000893009705F0000000c00000089000000890000008900000089", X"0000000c000000890000008937A7C5AC0000000c00000063000000890000008900000089", X"0000004900000089000000892B8CBCCC0000000d00000089000000890000008900000089", X"0000000e0000008900000089322BCC770000000d00000049000000890000008900000089",
 X"0000000d000000890000008937A7C5AC0000000d00000063000000890000008900000089", X"000000490000000d000000892EDBE6FE0000000e00000089000000890000008900000089", X"0000000f000000890000008931CE288E0000000e00000049000000890000008900000089", X"0000000e000000890000008937A7C5AC0000000e00000063000000890000008900000089", X"000000490000000e000000892EDBE6FE0000000f00000089000000890000008900000089", X"0000001000000089000000893189705F0000000f00000049000000890000008900000089",X"0000000f000000890000008937A7C5AC0000000f00000063000000890000008900000089", X"000000490000000f000000892EDBE6FE0000001000000089000000890000008900000089", X"0000001100000089000000893109705F0000001000000049000000890000008900000089", X"00000010000000890000008937A7C5AC0000001000000063000000890000008900000089",
 X"0000004900000010000000892EDBE6FE0000001100000089000000890000008900000089", X"00000011000000890000008937A7C5AC0000001100000063000000890000008900000089", X"00000011000000620000008931ABCC770000001200000089000000890000008900000089", X"0000001000000062000000893A83126E0000001200000089000000890000008900000089", X"0000000f000000620000008931ABCC770000001200000089000000890000008900000089", X"0000000e000000620000008931ABCC770000001200000089000000890000008900000089",X"0000000d000000620000008931ABCC770000001200000089000000890000008900000089", X"0000001c000000620000008931ABCC770000001200000089000000890000008900000089", X"0000001b000000620000008931ABCC770000001200000089000000890000008900000089", X"0000001a000000620000008931ABCC770000001200000089000000890000008900000089",  
 X"00000019000000620000008931ABCC770000001200000089000000890000008900000089", X"00000018000000620000008931ABCC770000001200000089000000890000008900000089", X"00000017000000620000008931ABCC770000001200000089000000890000008900000089", X"00000016000000620000008931ABCC770000001200000089000000890000008900000089", X"00000015000000620000008931ABCC770000001200000089000000890000008900000089", X"00000014000000620000008931ABCC770000001200000089000000890000008900000089",X"00000013000000620000008931ABCC770000001200000089000000890000008900000089", X"0000000c000000620000008931ABCC770000001200000089000000890000008900000089", X"0000000b000000620000008931ABCC770000001200000089000000890000008900000089", X"0000000a000000620000008931ABCC770000001200000089000000890000008900000089",
 X"00000009000000620000008931ABCC770000001200000089000000890000008900000089", X"00000008000000620000008931ABCC770000001200000089000000890000008900000089", X"00000007000000620000008931ABCC770000001200000089000000890000008900000089", X"00000006000000620000008931ABCC770000001200000089000000890000008900000089", X"00000005000000620000008931ABCC770000001200000089000000890000008900000089", X"00000004000000620000008931ABCC770000001200000089000000890000008900000089",X"00000003000000620000008931ABCC770000001200000089000000890000008900000089", X"0000006500000089000000892B8CBCCC0000001200000089000000890000008900000089", X"00000013000000890000008937A7C5AC0000001300000063000000890000008900000089", X"0000001400000089000000893189705F0000001300000065000000890000008900000089",
 X"0000006500000013000000892EDBE6FE0000001400000089000000890000008900000089", X"00000014000000890000008937A7C5AC0000001400000063000000890000008900000089", X"00000015000000890000008931CE288E0000001400000065000000890000008900000089", X"0000006500000014000000892EDBE6FE0000001500000089000000890000008900000089", X"00000015000000890000008937A7C5AC0000001500000063000000890000008900000089", X"0000001600000089000000893209705F0000001500000065000000890000008900000089",X"0000006500000015000000892EDBE6FE0000001600000089000000890000008900000089", X"00000016000000890000008937A7C5AC0000001600000063000000890000008900000089", X"000000170000008900000089322BCC770000001600000063000000890000008900000089", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",  
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001",
 X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001", X"0000000a00000012000000013A83126E0000000300000012000000120000000100000001");

begin 
 process (clk,en,we) 
 begin 
if en='1' then
  if (clk'event and clk = '1') then
 	  --if en='1' then
 	   	if (we = '1') then 
 			RAM(conv_integer(a)) <= di; 
 		else
		    do(31 downto 0)  <= RAM(conv_integer(a))(287 downto 256);
			 do0(31 downto 0) <= RAM(conv_integer(a))(255 downto 224);
		    do1(31 downto 0) <= RAM(conv_integer(a))(223 downto 192);
		    do2(31 downto 0) <= RAM(conv_integer(a))(191 downto 160);
 			 do3(31 downto 0) <= RAM(conv_integer(a))(159 downto 128);
			 do4(31 downto 0) <= RAM(conv_integer(a))(127 downto 96);
			 do5(31 downto 0) <= RAM(conv_integer(a))(95 downto 64);
			 do6(31 downto 0) <= RAM(conv_integer(a))(63 downto 32);
			 do7(31 downto 0) <= RAM(conv_integer(a))(31 downto 0);
 		end if;	  
 	end if; 
  end if;	
 end process; 


end Behavioral;


