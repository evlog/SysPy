----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:44:16 11/15/2011 
-- Design Name: 
-- Module Name:    speciescopyTableFRM2X_2 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity speciescopyTableFRM2X_2 is
port (clk : in std_logic; 
 	we  : in std_logic; 
 	en  : in std_logic;
 	--ssr : in std_logic;
 	a,a1,a2,a3 : in std_logic_vector(31 downto 0); 
 	di1,di2,di3,di4  : in std_logic_vector(31 downto 0); 
 	do,do1,do2,do3 : out std_logic_vector(31 downto 0));
end speciescopyTableFRM2X_2;

architecture Behavioral of speciescopyTableFRM2X_2 is

type ram_type1 is array(0 to 511) of std_logic_vector(31 downto 0);
signal RAM1:ram_type1:= 
(X"40a00000", X"40a00000", X"42be0000", X"00000000", X"00000000", X"00000000",X"00000000",X"3f800000", X"3f800000", X"00000000",  
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"42c80000",X"42c80000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"00000000", X"43200000",
 X"42D20000", X"4446C000", X"42480000", X"446D8000", X"43960000", X"43200000",X"40A00000",X"00000000", X"00000000", X"41A00000",
 X"00000000", X"41C80000", X"00000000", X"41C80000", X"00000000", X"41F00000",X"00000000",X"41F00000", X"00000000", X"42200000",
 X"41700000", X"42200000", X"41A00000", X"40000000", X"00000000", X"00000000",X"42C80000",X"00000000", X"42C80000", X"00000000",  
 X"42c80000", X"00000000", X"42C80000", X"00000000", X"42c80000", X"00000000",X"42C80000",X"43960000", X"42c80000", X"42c80000",
 X"43480000", X"00000000", X"44960000", X"42A00000", X"00000000", X"3f800000",X"40000000",X"41200000", X"43AF0000", X"45BB8000",
 X"45960000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"00000000", X"00000000",  
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"44BB8000", X"41200000",
 X"444BC000", X"40A00000", X"00000000", X"00000000", X"00000000", X"40A00000",X"41A00000",X"00000000", X"3f800000", X"3f800000",
 X"45B4C800", X"41200000", X"00000000", X"00000000", X"44BB8000", X"43FA0000",X"00000000",X"00000000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"453B8000",X"00000000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000");
 
 type ram_type2 is array(0 to 511) of std_logic_vector(31 downto 0);
signal RAM2:ram_type2:= 
(X"40a00000", X"40a00000", X"42be0000", X"00000000", X"00000000", X"00000000",X"00000000",X"3f800000", X"3f800000", X"00000000",  
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"42c80000",X"42c80000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"00000000", X"43200000",
 X"42D20000", X"4446C000", X"42480000", X"446D8000", X"43960000", X"43200000",X"40A00000",X"00000000", X"00000000", X"41A00000",
 X"00000000", X"41C80000", X"00000000", X"41C80000", X"00000000", X"41F00000",X"00000000",X"41F00000", X"00000000", X"42200000",
 X"41700000", X"42200000", X"41A00000", X"40000000", X"00000000", X"00000000",X"42C80000",X"00000000", X"42C80000", X"00000000",  
 X"42c80000", X"00000000", X"42C80000", X"00000000", X"42c80000", X"00000000",X"42C80000",X"43960000", X"42c80000", X"42c80000",
 X"43480000", X"00000000", X"44960000", X"42A00000", X"00000000", X"3f800000",X"40000000",X"41200000", X"43AF0000", X"45BB8000",
 X"45960000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"00000000", X"00000000",  
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"44BB8000", X"41200000",
 X"444BC000", X"40A00000", X"00000000", X"00000000", X"00000000", X"40A00000",X"41A00000",X"00000000", X"3f800000", X"3f800000",
 X"45B4C800", X"41200000", X"00000000", X"00000000", X"44BB8000", X"43FA0000",X"00000000",X"00000000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"453B8000",X"00000000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000");
 
 type ram_type3 is array(0 to 511) of std_logic_vector(31 downto 0);
signal RAM3:ram_type3:= 
(X"40a00000", X"40a00000", X"42be0000", X"00000000", X"00000000", X"00000000",X"00000000",X"3f800000", X"3f800000", X"00000000",  
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"42c80000",X"42c80000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"00000000", X"43200000",
 X"42D20000", X"4446C000", X"42480000", X"446D8000", X"43960000", X"43200000",X"40A00000",X"00000000", X"00000000", X"41A00000",
 X"00000000", X"41C80000", X"00000000", X"41C80000", X"00000000", X"41F00000",X"00000000",X"41F00000", X"00000000", X"42200000",
 X"41700000", X"42200000", X"41A00000", X"40000000", X"00000000", X"00000000",X"42C80000",X"00000000", X"42C80000", X"00000000",  
 X"42c80000", X"00000000", X"42C80000", X"00000000", X"42c80000", X"00000000",X"42C80000",X"43960000", X"42c80000", X"42c80000",
 X"43480000", X"00000000", X"44960000", X"42A00000", X"00000000", X"3f800000",X"40000000",X"41200000", X"43AF0000", X"45BB8000",
 X"45960000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"00000000", X"00000000",  
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"44BB8000", X"41200000",
 X"444BC000", X"40A00000", X"00000000", X"00000000", X"00000000", X"40A00000",X"41A00000",X"00000000", X"3f800000", X"3f800000",
 X"45B4C800", X"41200000", X"00000000", X"00000000", X"44BB8000", X"43FA0000",X"00000000",X"00000000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"453B8000",X"00000000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000");
 
 type ram_type4 is array(0 to 511) of std_logic_vector(31 downto 0);
signal RAM4:ram_type4:= 
(X"40a00000", X"40a00000", X"42be0000", X"00000000", X"00000000", X"00000000",X"00000000",X"3f800000", X"3f800000", X"00000000",  
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"42c80000",X"42c80000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"00000000", X"43200000",
 X"42D20000", X"4446C000", X"42480000", X"446D8000", X"43960000", X"43200000",X"40A00000",X"00000000", X"00000000", X"41A00000",
 X"00000000", X"41C80000", X"00000000", X"41C80000", X"00000000", X"41F00000",X"00000000",X"41F00000", X"00000000", X"42200000",
 X"41700000", X"42200000", X"41A00000", X"40000000", X"00000000", X"00000000",X"42C80000",X"00000000", X"42C80000", X"00000000",  
 X"42c80000", X"00000000", X"42C80000", X"00000000", X"42c80000", X"00000000",X"42C80000",X"43960000", X"42c80000", X"42c80000",
 X"43480000", X"00000000", X"44960000", X"42A00000", X"00000000", X"3f800000",X"40000000",X"41200000", X"43AF0000", X"45BB8000",
 X"45960000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"00000000", X"00000000",  
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"00000000",X"00000000", X"44BB8000", X"41200000",
 X"444BC000", X"40A00000", X"00000000", X"00000000", X"00000000", X"40A00000",X"41A00000",X"00000000", X"3f800000", X"3f800000",
 X"45B4C800", X"41200000", X"00000000", X"00000000", X"44BB8000", X"43FA0000",X"00000000",X"00000000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"453B8000",X"00000000", X"00000000", X"00000000",
 X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",  
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000", X"42C80000", X"00000000", X"00000000", X"42480000",X"42C80000",X"00000000", X"00000000", X"42480000",
 X"42480000", X"42480000");

begin 
 process (clk,en,we) 
begin 
if en='1' then
  if (clk'event and clk = '1') then
 	  --if en='1' then
 	   	if (we = '1') then 
 			RAM1(conv_integer(a)) <= di1; 
			RAM2(conv_integer(a1)) <= di2;
			RAM3(conv_integer(a2)) <= di3;
			RAM4(conv_integer(a3)) <= di4;
			
 		else
 			 do(31 downto 0)  <= RAM1(conv_integer(a));
			 do1(31 downto 0) <= RAM1(conv_integer(a1));
			 do2(31 downto 0) <= RAM1(conv_integer(a2));
			 do3(31 downto 0) <= RAM1(conv_integer(a3));
			 
			 			 
 		end if;	  
 	end if; 
  end if;	
 end process; 

end Behavioral;


