----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:43:47 01/11/2010 
-- Design Name: 
-- Module Name:    sin_comp - sin_comp_beh 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sin_comp is
    Port ( clk : in std_logic;
			  ang_in : in  std_logic_vector (9 downto 0);
           sin_out : out  std_logic_vector (17 downto 0));
	 attribute MULT_STYLE : string;
	 attribute MULT_STYLE of sin_comp : entity is "block";
	 attribute ROM_EXTRACT : string;
	 attribute ROM_EXTRACT of sin_comp : entity is "yes";
	 attribute ROM_STYLE : string;
	 attribute ROM_STYLE of sin_comp : entity is "block";
end sin_comp;

architecture sin_comp_beh of sin_comp is

--signal test: array (0 to 3) of std_logic_vector(3 downto 0);

type ROM_TYPE is array(0 to 2047)of std_logic_vector(17 downto 0);

constant sin_lut : ROM_TYPE := (
"000000000000000000", "000000000000110010", "000000000001100101", "000000000010010111", "000000000011001001", 
"000000000011111100", "000000000100101110", "000000000101100000", "000000000110010011", "000000000111000101", 
"000000000111110111", "000000001000101001", "000000001001011100", "000000001010001110", "000000001011000000", 
"000000001011110011", "000000001100100101", "000000001101010111", "000000001110001010", "000000001110111100", 
"000000001111101110", "000000010000100001", "000000010001010011", "000000010010000101", "000000010010110111", 
"000000010011101010", "000000010100011100", "000000010101001110", "000000010110000001", "000000010110110011", 
"000000010111100101", "000000011000011000", "000000011001001010", "000000011001111100", "000000011010101111", 
"000000011011100001", "000000011100010011", "000000011101000101", "000000011101111000", "000000011110101010", 
"000000011111011100", "000000100000001111", "000000100001000001", "000000100001110011", "000000100010100101", 
"000000100011011000", "000000100100001010", "000000100100111100", "000000100101101111", "000000100110100001", 
"000000100111010011", "000000101000000101", "000000101000111000", "000000101001101010", "000000101010011100", 
"000000101011001110", "000000101100000001", "000000101100110011", "000000101101100101", "000000101110011000", 
"000000101111001010", "000000101111111100", "000000110000101110", "000000110001100001", "000000110010010011", 
"000000110011000101", "000000110011110111", "000000110100101010", "000000110101011100", "000000110110001110", 
"000000110111000000", "000000110111110011", "000000111000100101", "000000111001010111", "000000111010001001", 
"000000111010111100", "000000111011101110", "000000111100100000", "000000111101010010", "000000111110000100", 
"000000111110110111", "000000111111101001", "000001000000011011", "000001000001001101", "000001000001111111", 
"000001000010110010", "000001000011100100", "000001000100010110", "000001000101001000", "000001000101111011", 
"000001000110101101", "000001000111011111", "000001001000010001", "000001001001000011", "000001001001110101", 
"000001001010101000", "000001001011011010", "000001001100001100", "000001001100111110", "000001001101110000", 
"000001001110100011", "000001001111010101", "000001010000000111", "000001010000111001", "000001010001101011", 
"000001010010011101", "000001010011001111", "000001010100000010", "000001010100110100", "000001010101100110", 
"000001010110011000", "000001010111001010", "000001010111111100", "000001011000101110", "000001011001100001", 
"000001011010010011", "000001011011000101", "000001011011110111", "000001011100101001", "000001011101011011", 
"000001011110001101", "000001011110111111", "000001011111110001", "000001100000100100", "000001100001010110", 
"000001100010001000", "000001100010111010", "000001100011101100", "000001100100011110", "000001100101010000", 
"000001100110000010", "000001100110110100", "000001100111100110", "000001101000011000", "000001101001001010", 
"000001101001111100", "000001101010101110", "000001101011100000", "000001101100010010", "000001101101000100", 
"000001101101110110", "000001101110101001", "000001101111011011", "000001110000001101", "000001110000111111", 
"000001110001110001", "000001110010100011", "000001110011010101", "000001110100000111", "000001110100111001", 
"000001110101101011", "000001110110011100", "000001110111001110", "000001111000000000", "000001111000110010", 
"000001111001100100", "000001111010010110", "000001111011001000", "000001111011111010", "000001111100101100", 
"000001111101011110", "000001111110010000", "000001111111000010", "000001111111110100", "000010000000100110", 
"000010000001011000", "000010000010001010", "000010000010111100", "000010000011101101", "000010000100011111", 
"000010000101010001", "000010000110000011", "000010000110110101", "000010000111100111", "000010001000011001", 
"000010001001001011", "000010001001111100", "000010001010101110", "000010001011100000", "000010001100010010", 
"000010001101000100", "000010001101110110", "000010001110100111", "000010001111011001", "000010010000001011", 
"000010010000111101", "000010010001101111", "000010010010100001", "000010010011010010", "000010010100000100", 
"000010010100110110", "000010010101101000", "000010010110011001", "000010010111001011", "000010010111111101", 
"000010011000101111", "000010011001100000", "000010011010010010", "000010011011000100", "000010011011110110", 
"000010011100100111", "000010011101011001", "000010011110001011", "000010011110111101", "000010011111101110", 
"000010100000100000", "000010100001010010", "000010100010000011", "000010100010110101", "000010100011100111", 
"000010100100011000", "000010100101001010", "000010100101111100", "000010100110101101", "000010100111011111", 
"000010101000010001", "000010101001000010", "000010101001110100", "000010101010100101", "000010101011010111", 
"000010101100001001", "000010101100111010", "000010101101101100", "000010101110011101", "000010101111001111", 
"000010110000000001", "000010110000110010", "000010110001100100", "000010110010010101", "000010110011000111", 
"000010110011111000", "000010110100101010", "000010110101011011", "000010110110001101", "000010110110111110", 
"000010110111110000", "000010111000100001", "000010111001010011", "000010111010000100", "000010111010110110", 
"000010111011100111", "000010111100011001", "000010111101001010", "000010111101111100", "000010111110101101", 
"000010111111011111", "000011000000010000", "000011000001000001", "000011000001110011", "000011000010100100", 
"000011000011010110", "000011000100000111", "000011000100111000", "000011000101101010", "000011000110011011", 
"000011000111001100", "000011000111111110", "000011001000101111", "000011001001100000", "000011001010010010", 
"000011001011000011", "000011001011110100", "000011001100100110", "000011001101010111", "000011001110001000", 
"000011001110111010", "000011001111101011", "000011010000011100", "000011010001001101", "000011010001111111", 
"000011010010110000", "000011010011100001", "000011010100010010", "000011010101000100", "000011010101110101", 
"000011010110100110", "000011010111010111", "000011011000001000", "000011011000111010", "000011011001101011", 
"000011011010011100", "000011011011001101", "000011011011111110", "000011011100101111", "000011011101100000", 
"000011011110010010", "000011011111000011", "000011011111110100", "000011100000100101", "000011100001010110", 
"000011100010000111", "000011100010111000", "000011100011101001", "000011100100011010", "000011100101001011", 
"000011100101111100", "000011100110101101", "000011100111011110", "000011101000001111", "000011101001000000", 
"000011101001110001", "000011101010100010", "000011101011010011", "000011101100000100", "000011101100110101", 
"000011101101100110", "000011101110010111", "000011101111001000", "000011101111111001", "000011110000101010", 
"000011110001011011", "000011110010001100", "000011110010111100", "000011110011101101", "000011110100011110", 
"000011110101001111", "000011110110000000", "000011110110110001", "000011110111100010", "000011111000010010", 
"000011111001000011", "000011111001110100", "000011111010100101", "000011111011010110", "000011111100000110", 
"000011111100110111", "000011111101101000", "000011111110011001", "000011111111001001", "000011111111111010", 
"000100000000101011", "000100000001011011", "000100000010001100", "000100000010111101", "000100000011101110", 
"000100000100011110", "000100000101001111", "000100000101111111", "000100000110110000", "000100000111100001", 
"000100001000010001", "000100001001000010", "000100001001110011", "000100001010100011", "000100001011010100", 
"000100001100000100", "000100001100110101", "000100001101100101", "000100001110010110", "000100001111000110", 
"000100001111110111", "000100010000100111", "000100010001011000", "000100010010001000", "000100010010111001", 
"000100010011101001", "000100010100011010", "000100010101001010", "000100010101111011", "000100010110101011", 
"000100010111011100", "000100011000001100", "000100011000111100", "000100011001101101", "000100011010011101", 
"000100011011001101", "000100011011111110", "000100011100101110", "000100011101011110", "000100011110001111", 
"000100011110111111", "000100011111101111", "000100100000100000", "000100100001010000", "000100100010000000", 
"000100100010110000", "000100100011100001", "000100100100010001", "000100100101000001", "000100100101110001", 
"000100100110100001", "000100100111010010", "000100101000000010", "000100101000110010", "000100101001100010", 
"000100101010010010", "000100101011000010", "000100101011110011", "000100101100100011", "000100101101010011", 
"000100101110000011", "000100101110110011", "000100101111100011", "000100110000010011", "000100110001000011", 
"000100110001110011", "000100110010100011", "000100110011010011", "000100110100000011", "000100110100110011", 
"000100110101100011", "000100110110010011", "000100110111000011", "000100110111110011", "000100111000100011", 
"000100111001010011", "000100111010000011", "000100111010110010", "000100111011100010", "000100111100010010", 
"000100111101000010", "000100111101110010", "000100111110100010", "000100111111010001", "000101000000000001", 
"000101000000110001", "000101000001100001", "000101000010010001", "000101000011000000", "000101000011110000", 
"000101000100100000", "000101000101010000", "000101000101111111", "000101000110101111", "000101000111011111", 
"000101001000001110", "000101001000111110", "000101001001101110", "000101001010011101", "000101001011001101", 
"000101001011111100", "000101001100101100", "000101001101011100", "000101001110001011", "000101001110111011", 
"000101001111101010", "000101010000011010", "000101010001001001", "000101010001111001", "000101010010101000", 
"000101010011011000", "000101010100000111", "000101010100110111", "000101010101100110", "000101010110010110", 
"000101010111000101", "000101010111110100", "000101011000100100", "000101011001010011", "000101011010000010", 
"000101011010110010", "000101011011100001", "000101011100010001", "000101011101000000", "000101011101101111", 
"000101011110011110", "000101011111001110", "000101011111111101", "000101100000101100", "000101100001011011", 
"000101100010001011", "000101100010111010", "000101100011101001", "000101100100011000", "000101100101000111", 
"000101100101110110", "000101100110100110", "000101100111010101", "000101101000000100", "000101101000110011", 
"000101101001100010", "000101101010010001", "000101101011000000", "000101101011101111", "000101101100011110", 
"000101101101001101", "000101101101111100", "000101101110101011", "000101101111011010", "000101110000001001", 
"000101110000111000", "000101110001100111", "000101110010010110", "000101110011000101", "000101110011110100", 
"000101110100100011", "000101110101010001", "000101110110000000", "000101110110101111", "000101110111011110", 
"000101111000001101", "000101111000111100", "000101111001101010", "000101111010011001", "000101111011001000", 
"000101111011110111", "000101111100100101", "000101111101010100", "000101111110000011", "000101111110110001", 
"000101111111100000", "000110000000001111", "000110000000111101", "000110000001101100", "000110000010011010", 
"000110000011001001", "000110000011111000", "000110000100100110", "000110000101010101", "000110000110000011", 
"000110000110110010", "000110000111100000", "000110001000001111", "000110001000111101", "000110001001101100", 
"000110001010011010", "000110001011001001", "000110001011110111", "000110001100100101", "000110001101010100", 
"000110001110000010", "000110001110110000", "000110001111011111", "000110010000001101", "000110010000111011", 
"000110010001101010", "000110010010011000", "000110010011000110", "000110010011110101", "000110010100100011", 
"000110010101010001", "000110010101111111", "000110010110101101", "000110010111011011", "000110011000001010", 
"000110011000111000", "000110011001100110", "000110011010010100", "000110011011000010", "000110011011110000", 
"000110011100011110", "000110011101001100", "000110011101111010", "000110011110101000", "000110011111010110", 
"000110100000000100", "000110100000110010", "000110100001100000", "000110100010001110", "000110100010111100", 
"000110100011101010", "000110100100011000", "000110100101000110", "000110100101110100", "000110100110100001", 
"000110100111001111", "000110100111111101", "000110101000101011", "000110101001011001", "000110101010000110", 
"000110101010110100", "000110101011100010", "000110101100010000", "000110101100111101", "000110101101101011", 
"000110101110011001", "000110101111000110", "000110101111110100", "000110110000100010", "000110110001001111", 
"000110110001111101", "000110110010101010", "000110110011011000", "000110110100000101", "000110110100110011", 
"000110110101100000", "000110110110001110", "000110110110111011", "000110110111101001", "000110111000010110", 
"000110111001000100", "000110111001110001", "000110111010011110", "000110111011001100", "000110111011111001", 
"000110111100100110", "000110111101010100", "000110111110000001", "000110111110101110", "000110111111011100", 
"000111000000001001", "000111000000110110", "000111000001100011", "000111000010010000", "000111000010111110", 
"000111000011101011", "000111000100011000", "000111000101000101", "000111000101110010", "000111000110011111", 
"000111000111001100", "000111000111111001", "000111001000100111", "000111001001010100", "000111001010000001", 
"000111001010101110", "000111001011011011", "000111001100000111", "000111001100110100", "000111001101100001", 
"000111001110001110", "000111001110111011", "000111001111101000", "000111010000010101", "000111010001000010", 
"000111010001101110", "000111010010011011", "000111010011001000", "000111010011110101", "000111010100100010", 
"000111010101001110", "000111010101111011", "000111010110101000", "000111010111010100", "000111011000000001", 
"000111011000101110", "000111011001011010", "000111011010000111", "000111011010110100", "000111011011100000", 
"000111011100001101", "000111011100111001", "000111011101100110", "000111011110010010", "000111011110111111", 
"000111011111101011", "000111100000011000", "000111100001000100", "000111100001110000", "000111100010011101", 
"000111100011001001", "000111100011110110", "000111100100100010", "000111100101001110", "000111100101111010", 
"000111100110100111", "000111100111010011", "000111100111111111", "000111101000101011", "000111101001011000", 
"000111101010000100", "000111101010110000", "000111101011011100", "000111101100001000", "000111101100110100", 
"000111101101100001", "000111101110001101", "000111101110111001", "000111101111100101", "000111110000010001", 
"000111110000111101", "000111110001101001", "000111110010010101", "000111110011000001", "000111110011101101", 
"000111110100011000", "000111110101000100", "000111110101110000", "000111110110011100", "000111110111001000", 
"000111110111110100", "000111111000100000", "000111111001001011", "000111111001110111", "000111111010100011", 
"000111111011001111", "000111111011111010", "000111111100100110", "000111111101010010", "000111111101111101", 
"000111111110101001", "000111111111010100", "001000000000000000", "001000000000101100", "001000000001010111", 
"001000000010000011", "001000000010101110", "001000000011011010", "001000000100000101", "001000000100110001", 
"001000000101011100", "001000000110000111", "001000000110110011", "001000000111011110", "001000001000001001", 
"001000001000110101", "001000001001100000", "001000001010001011", "001000001010110111", "001000001011100010", 
"001000001100001101", "001000001100111000", "001000001101100100", "001000001110001111", "001000001110111010", 
"001000001111100101", "001000010000010000", "001000010000111011", "001000010001100110", "001000010010010001", 
"001000010010111100", "001000010011100111", "001000010100010010", "001000010100111101", "001000010101101000", 
"001000010110010011", "001000010110111110", "001000010111101001", "001000011000010100", "001000011000111111", 
"001000011001101010", "001000011010010100", "001000011010111111", "001000011011101010", "001000011100010101", 
"001000011100111111", "001000011101101010", "001000011110010101", "001000011111000000", "001000011111101010", 
"001000100000010101", "001000100000111111", "001000100001101010", "001000100010010101", "001000100010111111", 
"001000100011101010", "001000100100010100", "001000100100111111", "001000100101101001", "001000100110010100", 
"001000100110111110", "001000100111101000", "001000101000010011", "001000101000111101", "001000101001100111", 
"001000101010010010", "001000101010111100", "001000101011100110", "001000101100010001", "001000101100111011", 
"001000101101100101", "001000101110001111", "001000101110111001", "001000101111100100", "001000110000001110", 
"001000110000111000", "001000110001100010", "001000110010001100", "001000110010110110", "001000110011100000", 
"001000110100001010", "001000110100110100", "001000110101011110", "001000110110001000", "001000110110110010", 
"001000110111011100", "001000111000000110", "001000111000101111", "001000111001011001", "001000111010000011", 
"001000111010101101", "001000111011010111", "001000111100000000", "001000111100101010", "001000111101010100", 
"001000111101111101", "001000111110100111", "001000111111010001", "001000111111111010", "001001000000100100", 
"001001000001001101", "001001000001110111", "001001000010100001", "001001000011001010", "001001000011110100", 
"001001000100011101", "001001000101000110", "001001000101110000", "001001000110011001", "001001000111000011", 
"001001000111101100", "001001001000010101", "001001001000111111", "001001001001101000", "001001001010010001", 
"001001001010111010", "001001001011100100", "001001001100001101", "001001001100110110", "001001001101011111", 
"001001001110001000", "001001001110110001", "001001001111011010", "001001010000000100", "001001010000101101", 
"001001010001010110", "001001010001111111", "001001010010101000", "001001010011010001", "001001010011111001", 
"001001010100100010", "001001010101001011", "001001010101110100", "001001010110011101", "001001010111000110", 
"001001010111101111", "001001011000010111", "001001011001000000", "001001011001101001", "001001011010010010", 
"001001011010111010", "001001011011100011", "001001011100001011", "001001011100110100", "001001011101011101", 
"001001011110000101", "001001011110101110", "001001011111010110", "001001011111111111", "001001100000100111", 
"001001100001010000", "001001100001111000", "001001100010100001", "001001100011001001", "001001100011110001", 
"001001100100011010", "001001100101000010", "001001100101101010", "001001100110010011", "001001100110111011", 
"001001100111100011", "001001101000001011", "001001101000110011", "001001101001011100", "001001101010000100", 
"001001101010101100", "001001101011010100", "001001101011111100", "001001101100100100", "001001101101001100", 
"001001101101110100", "001001101110011100", "001001101111000100", "001001101111101100", "001001110000010100", 
"001001110000111100", "001001110001100011", "001001110010001011", "001001110010110011", "001001110011011011", 
"001001110100000010", "001001110100101010", "001001110101010010", "001001110101111010", "001001110110100001", 
"001001110111001001", "001001110111110001", "001001111000011000", "001001111001000000", "001001111001100111", 
"001001111010001111", "001001111010110110", "001001111011011110", "001001111100000101", "001001111100101101", 
"001001111101010100", "001001111101111011", "001001111110100011", "001001111111001010", "001001111111110001", 
"001010000000011001", "001010000001000000", "001010000001100111", "001010000010001110", "001010000010110101", 
"001010000011011101", "001010000100000100", "001010000100101011", "001010000101010010", "001010000101111001", 
"001010000110100000", "001010000111000111", "001010000111101110", "001010001000010101", "001010001000111100", 
"001010001001100011", "001010001010001010", "001010001010110000", "001010001011010111", "001010001011111110", 
"001010001100100101", "001010001101001100", "001010001101110010", "001010001110011001", "001010001111000000", 
"001010001111100110", "001010010000001101", "001010010000110100", "001010010001011010", "001010010010000001", 
"001010010010100111", "001010010011001110", "001010010011110100", "001010010100011011", "001010010101000001", 
"001010010101101000", "001010010110001110", "001010010110110100", "001010010111011011", "001010011000000001", 
"001010011000100111", "001010011001001110", "001010011001110100", "001010011010011010", "001010011011000000", 
"001010011011100111", "001010011100001101", "001010011100110011", "001010011101011001", "001010011101111111", 
"001010011110100101", "001010011111001011", "001010011111110001", "001010100000010111", "001010100000111101", 
"001010100001100011", "001010100010001001", "001010100010101111", "001010100011010100", "001010100011111010", 
"001010100100100000", "001010100101000110", "001010100101101011", "001010100110010001", "001010100110110111", 
"001010100111011100", "001010101000000010", "001010101000101000", "001010101001001101", "001010101001110011", 
"001010101010011000", "001010101010111110", "001010101011100011", "001010101100001001", "001010101100101110", 
"001010101101010100", "001010101101111001", "001010101110011110", "001010101111000100", "001010101111101001", 
"001010110000001110", "001010110000110011", "001010110001011001", "001010110001111110", "001010110010100011", 
"001010110011001000", "001010110011101101", "001010110100010010", "001010110100110111", "001010110101011100", 
"001010110110000001", "001010110110100110", "001010110111001011", "001010110111110000", "001010111000010101", 
"001010111000111010", "001010111001011111", "001010111010000100", "001010111010101001", "001010111011001101", 
"001010111011110010", "001010111100010111", "001010111100111100", "001010111101100000", "001010111110000101", 
"001010111110101001", "001010111111001110", "001010111111110011", "001011000000010111", "001011000000111100", 
"001011000001100000", "001011000010000101", "001011000010101001", "001011000011001101", "001011000011110010", 
"001011000100010110", "001011000100111010", "001011000101011111", "001011000110000011", "001011000110100111", 
"001011000111001011", "001011000111110000", "001011001000010100", "001011001000111000", "001011001001011100", 
"001011001010000000", "001011001010100100", "001011001011001000", "001011001011101100", "001011001100010000", 
"001011001100110100", "001011001101011000", "001011001101111100", "001011001110100000", "001011001111000100", 
"001011001111100111", "001011010000001011", "001011010000101111", "001011010001010011", "001011010001110110", 
"001011010010011010", "001011010010111110", "001011010011100001", "001011010100000101", "001011010100101001", 
"001011010101001100", "001011010101110000", "001011010110010011", "001011010110110110", "001011010111011010", 
"001011010111111101", "001011011000100001", "001011011001000100", "001011011001100111", "001011011010001011", 
"001011011010101110", "001011011011010001", "001011011011110100", "001011011100011000", "001011011100111011", 
"001011011101011110", "001011011110000001", "001011011110100100", "001011011111000111", "001011011111101010", 
"001011100000001101", "001011100000110000", "001011100001010011", "001011100001110110", "001011100010011001", 
"001011100010111100", "001011100011011110", "001011100100000001", "001011100100100100", "001011100101000111", 
"001011100101101001", "001011100110001100", "001011100110101111", "001011100111010001", "001011100111110100", 
"001011101000010110", "001011101000111001", "001011101001011011", "001011101001111110", "001011101010100000", 
"001011101011000011", "001011101011100101", "001011101100001000", "001011101100101010", "001011101101001100", 
"001011101101101111", "001011101110010001", "001011101110110011", "001011101111010101", "001011101111110111", 
"001011110000011010", "001011110000111100", "001011110001011110", "001011110010000000", "001011110010100010", 
"001011110011000100", "001011110011100110", "001011110100001000", "001011110100101010", "001011110101001100", 
"001011110101101101", "001011110110001111", "001011110110110001", "001011110111010011", "001011110111110101", 
"001011111000010110", "001011111000111000", "001011111001011010", "001011111001111011", "001011111010011101", 
"001011111010111110", "001011111011100000", "001011111100000010", "001011111100100011", "001011111101000100", 
"001011111101100110", "001011111110000111", "001011111110101001", "001011111111001010", "001011111111101011", 
"001100000000001101", "001100000000101110", "001100000001001111", "001100000001110000", "001100000010010001", 
"001100000010110011", "001100000011010100", "001100000011110101", "001100000100010110", "001100000100110111", 
"001100000101011000", "001100000101111001", "001100000110011010", "001100000110111011", "001100000111011100", 
"001100000111111100", "001100001000011101", "001100001000111110", "001100001001011111", "001100001001111111", 
"001100001010100000", "001100001011000001", "001100001011100001", "001100001100000010", "001100001100100011", 
"001100001101000011", "001100001101100100", "001100001110000100", "001100001110100101", "001100001111000101", 
"001100001111100110", "001100010000000110", "001100010000100110", "001100010001000111", "001100010001100111", 
"001100010010000111", "001100010010100111", "001100010011001000", "001100010011101000", "001100010100001000", 
"001100010100101000", "001100010101001000", "001100010101101000", "001100010110001000", "001100010110101000", 
"001100010111001000", "001100010111101000", "001100011000001000", "001100011000101000", "001100011001001000", 
"001100011001100111", "001100011010000111", "001100011010100111", "001100011011000111", "001100011011100110", 
"001100011100000110", "001100011100100110", "001100011101000101", "001100011101100101", "001100011110000100", 
"001100011110100100", "001100011111000011", "001100011111100011", "001100100000000010", "001100100000100010", 
"001100100001000001", "001100100001100000", "001100100010000000", "001100100010011111", "001100100010111110", 
"001100100011011101", "001100100011111101", "001100100100011100", "001100100100111011", "001100100101011010", 
"001100100101111001", "001100100110011000", "001100100110110111", "001100100111010110", "001100100111110101", 
"001100101000010100", "001100101000110011", "001100101001010001", "001100101001110000", "001100101010001111", 
"001100101010101110", "001100101011001101", "001100101011101011", "001100101100001010", "001100101100101001", 
"001100101101000111", "001100101101100110", "001100101110000100", "001100101110100011", "001100101111000001", 
"001100101111100000", "001100101111111110", "001100110000011100", "001100110000111011", "001100110001011001", 
"001100110001110111", "001100110010010110", "001100110010110100", "001100110011010010", "001100110011110000", 
"001100110100001110", "001100110100101101", "001100110101001011", "001100110101101001", "001100110110000111", 
"001100110110100101", "001100110111000011", "001100110111100000", "001100110111111110", "001100111000011100", 
"001100111000111010", "001100111001011000", "001100111001110110", "001100111010010011", "001100111010110001", 
"001100111011001111", "001100111011101100", "001100111100001010", "001100111100101000", "001100111101000101", 
"001100111101100011", "001100111110000000", "001100111110011110", "001100111110111011", "001100111111011000", 
"001100111111110110", "001101000000010011", "001101000000110000", "001101000001001110", "001101000001101011", 
"001101000010001000", "001101000010100101", "001101000011000010", "001101000011011111", "001101000011111101", 
"001101000100011010", "001101000100110111", "001101000101010100", "001101000101110001", "001101000110001101", 
"001101000110101010", "001101000111000111", "001101000111100100", "001101001000000001", "001101001000011110", 
"001101001000111010", "001101001001010111", "001101001001110100", "001101001010010000", "001101001010101101", 
"001101001011001001", "001101001011100110", "001101001100000010", "001101001100011111", "001101001100111011", 
"001101001101011000", "001101001101110100", "001101001110010001", "001101001110101101", "001101001111001001", 
"001101001111100101", "001101010000000010", "001101010000011110", "001101010000111010", "001101010001010110", 
"001101010001110010", "001101010010001110", "001101010010101010", "001101010011000110", "001101010011100010", 
"001101010011111110", "001101010100011010", "001101010100110110", "001101010101010010", "001101010101101101", 
"001101010110001001", "001101010110100101", "001101010111000001", "001101010111011100", "001101010111111000", 
"001101011000010100", "001101011000101111", "001101011001001011", "001101011001100110", "001101011010000010", 
"001101011010011101", "001101011010111001", "001101011011010100", "001101011011101111", "001101011100001011", 
"001101011100100110", "001101011101000001", "001101011101011100", "001101011101111000", "001101011110010011", 
"001101011110101110", "001101011111001001", "001101011111100100", "001101011111111111", "001101100000011010", 
"001101100000110101", "001101100001010000", "001101100001101011", "001101100010000110", "001101100010100000", 
"001101100010111011", "001101100011010110", "001101100011110001", "001101100100001011", "001101100100100110", 
"001101100101000001", "001101100101011011", "001101100101110110", "001101100110010000", "001101100110101011", 
"001101100111000101", "001101100111100000", "001101100111111010", "001101101000010101", "001101101000101111", 
"001101101001001001", "001101101001100100", "001101101001111110", "001101101010011000", "001101101010110010", 
"001101101011001100", "001101101011100110", "001101101100000000", "001101101100011010", "001101101100110100", 
"001101101101001110", "001101101101101000", "001101101110000010", "001101101110011100", "001101101110110110", 
"001101101111010000", "001101101111101010", "001101110000000011", "001101110000011101", "001101110000110111", 
"001101110001010000", "001101110001101010", "001101110010000100", "001101110010011101", "001101110010110111", 
"001101110011010000", "001101110011101010", "001101110100000011", "001101110100011100", "001101110100110110", 
"001101110101001111", "001101110101101000", "001101110110000001", "001101110110011011", "001101110110110100", 
"001101110111001101", "001101110111100110", "001101110111111111", "001101111000011000", "001101111000110001", 
"001101111001001010", "001101111001100011", "001101111001111100", "001101111010010101", "001101111010101110", 
"001101111011000111", "001101111011011111", "001101111011111000", "001101111100010001", "001101111100101001", 
"001101111101000010", "001101111101011011", "001101111101110011", "001101111110001100", "001101111110100100", 
"001101111110111101", "001101111111010101", "001101111111101110", "001110000000000110", "001110000000011110", 
"001110000000110111", "001110000001001111", "001110000001100111", "001110000001111111", "001110000010010111", 
"001110000010110000", "001110000011001000", "001110000011100000", "001110000011111000", "001110000100010000", 
"001110000100101000", "001110000101000000", "001110000101011000", "001110000101101111", "001110000110000111", 
"001110000110011111", "001110000110110111", "001110000111001110", "001110000111100110", "001110000111111110", 
"001110001000010101", "001110001000101101", "001110001001000101", "001110001001011100", "001110001001110100", 
"001110001010001011", "001110001010100010", "001110001010111010", "001110001011010001", "001110001011101000", 
"001110001100000000", "001110001100010111", "001110001100101110", "001110001101000101", "001110001101011101", 
"001110001101110100", "001110001110001011", "001110001110100010", "001110001110111001", "001110001111010000", 
"001110001111100111", "001110001111111110", "001110010000010100", "001110010000101011", "001110010001000010", 
"001110010001011001", "001110010001110000", "001110010010000110", "001110010010011101", "001110010010110100", 
"001110010011001010", "001110010011100001", "001110010011110111", "001110010100001110", "001110010100100100", 
"001110010100111011", "001110010101010001", "001110010101100111", "001110010101111110", "001110010110010100", 
"001110010110101010", "001110010111000000", "001110010111010111", "001110010111101101", "001110011000000011", 
"001110011000011001", "001110011000101111", "001110011001000101", "001110011001011011", "001110011001110001", 
"001110011010000111", "001110011010011101", "001110011010110010", "001110011011001000", "001110011011011110", 
"001110011011110100", "001110011100001001", "001110011100011111", "001110011100110101", "001110011101001010", 
"001110011101100000", "001110011101110101", "001110011110001011", "001110011110100000", "001110011110110110", 
"001110011111001011", "001110011111100000", "001110011111110110", "001110100000001011", "001110100000100000", 
"001110100000110101", "001110100001001010", "001110100001100000", "001110100001110101", "001110100010001010", 
"001110100010011111", "001110100010110100", "001110100011001001", "001110100011011110", "001110100011110011", 
"001110100100000111", "001110100100011100", "001110100100110001", "001110100101000110", "001110100101011010", 
"001110100101101111", "001110100110000100", "001110100110011000", "001110100110101101", "001110100111000001", 
"001110100111010110", "001110100111101010", "001110100111111111", "001110101000010011", "001110101000101000", 
"001110101000111100", "001110101001010000", "001110101001100100", "001110101001111001", "001110101010001101", 
"001110101010100001", "001110101010110101", "001110101011001001", "001110101011011101", "001110101011110001", 
"001110101100000101", "001110101100011001", "001110101100101101", "001110101101000001", "001110101101010101", 
"001110101101101000", "001110101101111100", "001110101110010000", "001110101110100100", "001110101110110111", 
"001110101111001011", "001110101111011110", "001110101111110010", "001110110000000101", "001110110000011001", 
"001110110000101100", "001110110001000000", "001110110001010011", "001110110001100110", "001110110001111010", 
"001110110010001101", "001110110010100000", "001110110010110011", "001110110011000111", "001110110011011010", 
"001110110011101101", "001110110100000000", "001110110100010011", "001110110100100110", "001110110100111001", 
"001110110101001100", "001110110101011110", "001110110101110001", "001110110110000100", "001110110110010111", 
"001110110110101010", "001110110110111100", "001110110111001111", "001110110111100001", "001110110111110100", 
"001110111000000111", "001110111000011001", "001110111000101100", "001110111000111110", "001110111001010000", 
"001110111001100011", "001110111001110101", "001110111010000111", "001110111010011010", "001110111010101100", 
"001110111010111110", "001110111011010000", "001110111011100010", "001110111011110100", "001110111100000110", 
"001110111100011000", "001110111100101010", "001110111100111100", "001110111101001110", "001110111101100000", 
"001110111101110010", "001110111110000100", "001110111110010101", "001110111110100111", "001110111110111001", 
"001110111111001010", "001110111111011100", "001110111111101101", "001110111111111111", "001111000000010001", 
"001111000000100010", "001111000000110011", "001111000001000101", "001111000001010110", "001111000001100111", 
"001111000001111001", "001111000010001010", "001111000010011011", "001111000010101100", "001111000010111101", 
"001111000011001111", "001111000011100000", "001111000011110001", "001111000100000010", "001111000100010011", 
"001111000100100011", "001111000100110100", "001111000101000101", "001111000101010110", "001111000101100111", 
"001111000101110111", "001111000110001000", "001111000110011001", "001111000110101001", "001111000110111010", 
"001111000111001011", "001111000111011011", "001111000111101100", "001111000111111100", "001111001000001100", 
"001111001000011101", "001111001000101101", "001111001000111101", "001111001001001110", "001111001001011110", 
"001111001001101110", "001111001001111110", "001111001010001110", "001111001010011110", "001111001010101110", 
"001111001010111110", "001111001011001110", "001111001011011110", "001111001011101110", "001111001011111110", 
"001111001100001110", "001111001100011110", "001111001100101101", "001111001100111101", "001111001101001101", 
"001111001101011100", "001111001101101100", "001111001101111100", "001111001110001011", "001111001110011011", 
"001111001110101010", "001111001110111001", "001111001111001001", "001111001111011000", "001111001111100111", 
"001111001111110111", "001111010000000110", "001111010000010101", "001111010000100100", "001111010000110011", 
"001111010001000010", "001111010001010010", "001111010001100001", "001111010001101111", "001111010001111110", 
"001111010010001101", "001111010010011100", "001111010010101011", "001111010010111010", "001111010011001001", 
"001111010011010111", "001111010011100110", "001111010011110101", "001111010100000011", "001111010100010010", 
"001111010100100000", "001111010100101111", "001111010100111101", "001111010101001100", "001111010101011010", 
"001111010101101000", "001111010101110111", "001111010110000101", "001111010110010011", "001111010110100001", 
"001111010110101111", "001111010110111110", "001111010111001100", "001111010111011010", "001111010111101000", 
"001111010111110110", "001111011000000100", "001111011000010010", "001111011000011111", "001111011000101101", 
"001111011000111011", "001111011001001001", "001111011001010110", "001111011001100100", "001111011001110010", 
"001111011001111111", "001111011010001101", "001111011010011010", "001111011010101000", "001111011010110101", 
"001111011011000011", "001111011011010000", "001111011011011110", "001111011011101011", "001111011011111000", 
"001111011100000101", "001111011100010011", "001111011100100000", "001111011100101101", "001111011100111010", 
"001111011101000111", "001111011101010100", "001111011101100001", "001111011101101110", "001111011101111011", 
"001111011110001000", "001111011110010100", "001111011110100001", "001111011110101110", "001111011110111011", 
"001111011111000111", "001111011111010100", "001111011111100000", "001111011111101101", "001111011111111010", 
"001111100000000110", "001111100000010010", "001111100000011111", "001111100000101011", "001111100000111000", 
"001111100001000100", "001111100001010000", "001111100001011100", "001111100001101001", "001111100001110101", 
"001111100010000001", "001111100010001101", "001111100010011001", "001111100010100101", "001111100010110001", 
"001111100010111101", "001111100011001001", "001111100011010100", "001111100011100000", "001111100011101100", 
"001111100011111000", "001111100100000011", "001111100100001111", "001111100100011011", "001111100100100110", 
"001111100100110010", "001111100100111101", "001111100101001001", "001111100101010100", "001111100101100000", 
"001111100101101011", "001111100101110110", "001111100110000010", "001111100110001101", "001111100110011000", 
"001111100110100011", "001111100110101110", "001111100110111001", "001111100111000101", "001111100111010000", 
"001111100111011011", "001111100111100101", "001111100111110000", "001111100111111011", "001111101000000110", 
"001111101000010001", "001111101000011100", "001111101000100110", "001111101000110001", "001111101000111100", 
"001111101001000110", "001111101001010001", "001111101001011011", "001111101001100110", "001111101001110000", 
"001111101001111011", "001111101010000101", "001111101010001111", "001111101010011010", "001111101010100100", 
"001111101010101110", "001111101010111000", "001111101011000010", "001111101011001101", "001111101011010111", 
"001111101011100001", "001111101011101011", "001111101011110101", "001111101011111111", "001111101100001000", 
"001111101100010010", "001111101100011100", "001111101100100110", "001111101100110000", "001111101100111001", 
"001111101101000011", "001111101101001101", "001111101101010110", "001111101101100000", "001111101101101001", 
"001111101101110011", "001111101101111100", "001111101110000101", "001111101110001111", "001111101110011000", 
"001111101110100001", "001111101110101011", "001111101110110100", "001111101110111101", "001111101111000110", 
"001111101111001111", "001111101111011000", "001111101111100001", "001111101111101010", "001111101111110011", 
"001111101111111100", "001111110000000101", "001111110000001110", "001111110000010111", "001111110000011111", 
"001111110000101000", "001111110000110001", "001111110000111001", "001111110001000010", "001111110001001010", 
"001111110001010011", "001111110001011011", "001111110001100100", "001111110001101100", "001111110001110101", 
"001111110001111101", "001111110010000101", "001111110010001101", "001111110010010110", "001111110010011110", 
"001111110010100110", "001111110010101110", "001111110010110110", "001111110010111110", "001111110011000110", 
"001111110011001110", "001111110011010110", "001111110011011110", "001111110011100110", "001111110011101101", 
"001111110011110101", "001111110011111101", "001111110100000101", "001111110100001100", "001111110100010100", 
"001111110100011011", "001111110100100011", "001111110100101010", "001111110100110010", "001111110100111001", 
"001111110101000001", "001111110101001000", "001111110101001111", "001111110101010111", "001111110101011110", 
"001111110101100101", "001111110101101100", "001111110101110011", "001111110101111010", "001111110110000001", 
"001111110110001000", "001111110110001111", "001111110110010110", "001111110110011101", "001111110110100100", 
"001111110110101011", "001111110110110001", "001111110110111000", "001111110110111111", "001111110111000101", 
"001111110111001100", "001111110111010011", "001111110111011001", "001111110111100000", "001111110111100110", 
"001111110111101100", "001111110111110011", "001111110111111001", "001111111000000000", "001111111000000110", 
"001111111000001100", "001111111000010010", "001111111000011000", "001111111000011110", "001111111000100100", 
"001111111000101011", "001111111000110001", "001111111000110110", "001111111000111100", "001111111001000010", 
"001111111001001000", "001111111001001110", "001111111001010100", "001111111001011001", "001111111001011111", 
"001111111001100101", "001111111001101010", "001111111001110000", "001111111001110101", "001111111001111011", 
"001111111010000000", "001111111010000110", "001111111010001011", "001111111010010001", "001111111010010110", 
"001111111010011011", "001111111010100000", "001111111010100101", "001111111010101011", "001111111010110000", 
"001111111010110101", "001111111010111010", "001111111010111111", "001111111011000100", "001111111011001001", 
"001111111011001110", "001111111011010010", "001111111011010111", "001111111011011100", "001111111011100001", 
"001111111011100101", "001111111011101010", "001111111011101111", "001111111011110011", "001111111011111000", 
"001111111011111100", "001111111100000001", "001111111100000101", "001111111100001010", "001111111100001110", 
"001111111100010010", "001111111100010110", "001111111100011011", "001111111100011111", "001111111100100011", 
"001111111100100111", "001111111100101011", "001111111100101111", "001111111100110011", "001111111100110111", 
"001111111100111011", "001111111100111111", "001111111101000011", "001111111101000111", "001111111101001010", 
"001111111101001110", "001111111101010010", "001111111101010101", "001111111101011001", "001111111101011101", 
"001111111101100000", "001111111101100100", "001111111101100111", "001111111101101010", "001111111101101110", 
"001111111101110001", "001111111101110101", "001111111101111000", "001111111101111011", "001111111101111110", 
"001111111110000001", "001111111110000100", "001111111110000111", "001111111110001011", "001111111110001110", 
"001111111110010000", "001111111110010011", "001111111110010110", "001111111110011001", "001111111110011100", 
"001111111110011111", "001111111110100001", "001111111110100100", "001111111110100111", "001111111110101001", 
"001111111110101100", "001111111110101110", "001111111110110001", "001111111110110011", "001111111110110110", 
"001111111110111000", "001111111110111010", "001111111110111101", "001111111110111111", "001111111111000001", 
"001111111111000011", "001111111111000110", "001111111111001000", "001111111111001010", "001111111111001100", 
"001111111111001110", "001111111111010000", "001111111111010010", "001111111111010100", "001111111111010101", 
"001111111111010111", "001111111111011001", "001111111111011011", "001111111111011100", "001111111111011110", 
"001111111111100000", "001111111111100001", "001111111111100011", "001111111111100100", "001111111111100110", 
"001111111111100111", "001111111111101000", "001111111111101010", "001111111111101011", "001111111111101100", 
"001111111111101101", "001111111111101111", "001111111111110000", "001111111111110001", "001111111111110010", 
"001111111111110011", "001111111111110100", "001111111111110101", "001111111111110110", "001111111111110111", 
"001111111111110111", "001111111111111000", "001111111111111001", "001111111111111010", "001111111111111010", 
"001111111111111010", "001111111111111011", "001111111111111100", "001111111111111100", "001111111111111101", 
"001111111111111101", "001111111111111110", "001111111111111110", "001111111111111110", "001111111111111111", 
"001111111111111111", "001111111111111111", "001111111111111111", "001111111111111111", "001111111111111111",
"001111111111111111", "001111111111111111", "010000000000000000"); 

constant pi2 : std_logic_vector(9 downto 0) := "0001100101";
constant pi22 : std_logic_vector(9 downto 0) := "0011001001";
constant pi23 : std_logic_vector(9 downto 0) := "0100101110";
constant pi24 : std_logic_vector(9 downto 0) := "0110010010"; 
constant pi124 : std_logic_vector(9 downto 0) := "0000001010";

--signal sin_out_int : integer range 0 to 255;
signal ang_int : std_logic_vector(17 downto 0);
signal ang_in_int, temp1, temp3 : std_logic_vector(9 downto 0);
signal index0, index1, index2, sin_out_int, sin_out_int_neg : std_logic_vector(17 downto 0);
signal temp0, temp2 : std_logic_vector(19 downto 0);

begin

index0 <= (pi22 - ang_in_int) * "0001010001" + "0000000100";
index1 <= (ang_in_int - pi22) * "0001010001" + "0000000100";
index2 <= (pi24 - ang_in_int) * "0001010001" + "0000001000";

temp0 <= ang_in * pi124;
temp1 <= "00" & temp0(19 downto 12);
temp2 <= temp1 * pi24;
temp3 <= ang_in - temp2(9 downto 0);

ang_in_int <= ang_in when (ang_in <= pi24) else
              temp3;
				  

--ang_int <= ang_in_int * "000010100" + "000000100";

process(clk) begin
  if rising_edge(clk) then
  --if ((ang_in_int >= "000000000") and (ang_in_int < pi2)) then
	  if ang_in_int = "0000000000" then
			sin_out_int <= (others => '0');
			sin_out_int_neg <= (others => '0');
	  elsif ang_in_int /= "0000000000" then
			sin_out_int <= sin_lut(conv_integer(ang_int(10 downto 0)));
			sin_out_int_neg <= "000000000000000000" - sin_lut(conv_integer(ang_int(10 downto 0)));
	  end if;
  --elsif ((ang_in_int >= pi2) and (ang_in_int < pi22)) then
	--	sin_out <= sin_lut(conv_integer(index0(10 downto 0)));
  --elsif ((ang_in_int >= pi22) and (ang_in_int < pi23)) then
	--	sin_out <= ("000000000000000000" - sin_lut(conv_integer(index1(10 downto 0))));
  --elsif ((ang_in_int >= pi23) and (ang_in_int <= pi24)) then
--		sin_out <= ("000000000000000000" - sin_lut(conv_integer(index2(10 downto 0))));
  --else
	--	sin_out <= (others => '0');
  --end if;
  end if;
end process;

sin_out <= sin_out_int when ((ang_in_int >= "0000000000") and (ang_in_int < pi2)) else
			  sin_out_int when ((ang_in_int >= pi2) and (ang_in_int < pi22)) else
			  sin_out_int_neg when ((ang_in_int >= pi22) and (ang_in_int < pi23)) else
           sin_out_int_neg when ((ang_in_int >= pi23) and (ang_in_int <= pi24)) else
			  (others => '0');

ang_int <= (ang_in_int * "0001010001" + "0000000100") when ((ang_in_int >= "0000000000") and (ang_in_int < pi2)) else
			  index0 when ((ang_in_int >= pi2) and (ang_in_int < pi22)) else
			  index1 when ((ang_in_int >= pi22) and (ang_in_int < pi23)) else
           index2 when ((ang_in_int >= pi23) and (ang_in_int <= pi24)) else
			  (others => '0');

end sin_comp_beh;

