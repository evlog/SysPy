----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:12:53 09/13/2011 
-- Design Name: 
-- Module Name:    LOTKA_VOLTERA_STOICHIO - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LOTKA_VOLTERA_STOICHIO is
port (clk : in std_logic; 
 	we  : in std_logic; 
 	en  : in std_logic;
 	--ssr : in std_logic;
 	a   : in std_logic_vector(8 downto 0); 
 	di  : in std_logic_vector(255 downto 0); 
 	do0,do1,do2,do3,do4,do5,do6,do7  : out std_logic_vector(31 downto 0));
end LOTKA_VOLTERA_STOICHIO;

architecture Behavioral of LOTKA_VOLTERA_STOICHIO is

type ram_type is array(0 to 511) of std_logic_vector(255 downto 0);
signal RAM:ram_type:=
(X"3f80000000000000000000000000000000000000000000000000000000000000",X"bf8000003f800000000000000000000000000000000000000000000000000000", X"bf80000000000000000000000000000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"0000000000000000000000003f80000000000000000000000000000000000000", X"bf80000000000000000000003f8000003f800000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"000000000000000000000000000000003f800000000000000000000000000000",X"bf80000000000000000000003f8000003f800000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000", 
 X"000000000000000000000000000000003f800000000000000000000000000000",X"bf80000000000000000000003f8000003f800000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"0000000000000000000000003f80000000000000000000000000000000000000",X"c000000000000000000000003f80000000000000000000000000000000000000", X"000000000000000000000000000000003f800000000000000000000000000000",X"bf80000000000000000000003f8000003f800000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"000000000000000000000000000000003f800000000000000000000000000000", X"bf80000000000000000000003f8000003f800000000000000000000000000000",
 X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"0000000000000000000000003f80000000000000000000000000000000000000", X"bf80000000000000000000003f8000003f800000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"000000000000000000000000000000003f800000000000000000000000000000", X"bf80000000000000000000003f8000003f800000000000000000000000000000",X"bf800000bf800000000000003f8000003f800000000000000000000000000000",X"000000000000000000000000000000003f800000000000000000000000000000",X"c000000000000000000000003f80000000000000000000000000000000000000", X"bf80000000000000000000003f8000003f800000000000000000000000000000", 
 X"000000000000000000000000000000003f800000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"0000000000000000000000003f8000003f800000000000000000000000000000", X"000000000000000000000000000000003f800000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf80000000000000000000003f8000003f800000000000000000000000000000",X"0000000000000000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf80000000000000000000003f8000003f800000000000000000000000000000", X"000000000000000000000000000000003f800000000000000000000000000000",
 X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"0000000000000000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000",
 X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000", 
 X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"c000000000000000000000003f80000000000000000000000000000000000000",X"000000000000000000000000000000003f800000000000000000000000000000", X"bf80000000000000000000003f8000003f800000000000000000000000000000",
 X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"000000000000000000000000000000003f800000000000000000000000000000", X"bf80000000000000000000003f8000003f800000000000000000000000000000", X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"000000000000000000000000000000003f800000000000000000000000000000", X"bf80000000000000000000003f8000003f800000000000000000000000000000",X"bf800000bf800000000000003f80000000000000000000000000000000000000",X"000000000000000000000000000000003f800000000000000000000000000000",X"bf8000000000000000000000000000003f8000003f8000000000000000000000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", 
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", 
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", 
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", 
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", 
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", 
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", 
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", 
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", 
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", 
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000", X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",
 X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000",X"bf8000000000000000000000000000003f8000003f8000003f8000003f800000");

 begin 
 process (clk,en,we) 
 begin 
if en='1' then
  if (clk'event and clk = '1') then
 	  --if en='1' then
 	   	if (we = '1') then 
 			RAM(conv_integer(a)) <= di; 
 		else
		    do0(31 downto 0) <= RAM(conv_integer(a))(255 downto 224);
		    do1(31 downto 0) <= RAM(conv_integer(a))(223 downto 192);
		    do2(31 downto 0) <= RAM(conv_integer(a))(191 downto 160);
		    do3(31 downto 0) <= RAM(conv_integer(a))(159 downto 128);
 			 do4(31 downto 0) <= RAM(conv_integer(a))(127 downto 96);
			 do5(31 downto 0) <= RAM(conv_integer(a))(95 downto 64);
			 do6(31 downto 0) <= RAM(conv_integer(a))(63 downto 32);
			 do7(31 downto 0) <= RAM(conv_integer(a))(31 downto 0);
 		end if;	  
 	end if; 
  end if;	
 end process; 
end Behavioral;

